module Project_2_top (button, Clk, led, seg_sec, seg_tsec, seg_hsec);
	input [1:0] button;
	input Clk;
	output led;
	output [7:0] seg_sec;
	output [6:0] seg_tsec, seg_hsec;
	
endmodule 
